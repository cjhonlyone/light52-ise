--------------------------------------------------------------------------------
-- obj_code_pkg.vhdl -- Application object code in vhdl constant string format.
--------------------------------------------------------------------------------
-- Written by build_rom.py for project 'Blinker'.
--------------------------------------------------------------------------------
-- Copyright (C) 2012 Jose A. Ruiz
--
-- This source file may be used and distributed without
-- restriction provided that this copyright statement is not
-- removed from the file and that any derivative work contains
-- the original copyright notice and the associated disclaimer.
--
-- This source file is free software; you can redistribute it
-- and/or modify it under the terms of the GNU Lesser General
-- Public License as published by the Free Software Foundation;
-- either version 2.1 of the License, or (at your option) any
-- later version.
--
-- This source is distributed in the hope that it will be
-- useful, but WITHOUT ANY WARRANTY; without even the implied
-- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR
-- PURPOSE.  See the GNU Lesser General Public License for more
-- details.
--
-- You should have received a copy of the GNU Lesser General
-- Public License along with this source; if not, download it
-- from http://www.opencores.org/lgpl.shtml
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.light52_pkg.all;

package obj_code_pkg is

-- Size of XCODE memory in bytes.
constant XCODE_SIZE : natural := 8192;
-- Size of XDATA memory in bytes.
constant XDATA_SIZE : natural := 0;

-- Object code initialization constant.
constant object_code : t_obj_code(0 to 5684) := (
    X"02", X"00", X"3f", X"32", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"02", X"09", X"7f", X"02", X"00", 
    X"c2", X"e5", X"81", X"24", X"fc", X"c3", X"c8", X"c0", 
    X"e0", X"c0", X"82", X"e6", X"08", X"46", X"70", X"06", 
    X"e5", X"82", X"45", X"83", X"60", X"12", X"18", X"e5", 
    X"82", X"96", X"f5", X"82", X"08", X"e5", X"83", X"96", 
    X"42", X"82", X"08", X"e5", X"f0", X"96", X"45", X"82", 
    X"d0", X"82", X"c8", X"d0", X"e0", X"c8", X"22", X"75", 
    X"81", X"7c", X"12", X"14", X"f5", X"e5", X"82", X"60", 
    X"03", X"02", X"00", X"0e", X"79", X"00", X"e9", X"44", 
    X"00", X"60", X"1b", X"7a", X"00", X"90", X"16", X"35", 
    X"78", X"01", X"75", X"a0", X"00", X"e4", X"93", X"f2", 
    X"a3", X"08", X"b8", X"00", X"02", X"05", X"a0", X"d9", 
    X"f4", X"da", X"f2", X"75", X"a0", X"ff", X"e4", X"78", 
    X"ff", X"f6", X"d8", X"fd", X"78", X"00", X"e8", X"44", 
    X"00", X"60", X"0a", X"79", X"01", X"75", X"a0", X"00", 
    X"e4", X"f3", X"09", X"d8", X"fc", X"78", X"00", X"e8", 
    X"44", X"00", X"60", X"0c", X"79", X"00", X"90", X"00", 
    X"01", X"e4", X"f0", X"a3", X"d8", X"fc", X"d9", X"fa", 
    X"75", X"09", X"fc", X"75", X"0a", X"60", X"75", X"0b", 
    X"da", X"75", X"0c", X"f2", X"75", X"0d", X"66", X"75", 
    X"0e", X"b6", X"75", X"0f", X"be", X"75", X"10", X"e0", 
    X"75", X"11", X"fe", X"75", X"12", X"f6", X"75", X"13", 
    X"01", X"75", X"14", X"00", X"75", X"3b", X"00", X"02", 
    X"00", X"0e", X"12", X"08", X"a3", X"e4", X"f5", X"25", 
    X"f5", X"26", X"7b", X"15", X"7c", X"00", X"7d", X"40", 
    X"c0", X"05", X"c0", X"04", X"c0", X"03", X"74", X"f9", 
    X"c0", X"e0", X"74", X"14", X"c0", X"e0", X"74", X"80", 
    X"c0", X"e0", X"12", X"0c", X"13", X"15", X"81", X"15", 
    X"81", X"15", X"81", X"74", X"fb", X"c0", X"e0", X"74", 
    X"14", X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", 
    X"0c", X"13", X"15", X"81", X"15", X"81", X"15", X"81", 
    X"74", X"1e", X"c0", X"e0", X"74", X"15", X"c0", X"e0", 
    X"74", X"80", X"c0", X"e0", X"12", X"0c", X"13", X"15", 
    X"81", X"15", X"81", X"15", X"81", X"74", X"4a", X"c0", 
    X"e0", X"74", X"15", X"c0", X"e0", X"74", X"80", X"c0", 
    X"e0", X"12", X"0c", X"13", X"15", X"81", X"15", X"81", 
    X"15", X"81", X"d0", X"03", X"d0", X"04", X"d0", X"05", 
    X"20", X"9d", X"03", X"02", X"05", X"b4", X"aa", X"99", 
    X"7f", X"00", X"c0", X"07", X"c0", X"05", X"c0", X"04", 
    X"c0", X"03", X"c0", X"02", X"c0", X"25", X"c0", X"26", 
    X"c0", X"02", X"c0", X"07", X"74", X"7d", X"c0", X"e0", 
    X"74", X"15", X"c0", X"e0", X"74", X"80", X"c0", X"e0", 
    X"12", X"0c", X"13", X"e5", X"81", X"24", X"f9", X"f5", 
    X"81", X"d0", X"02", X"d0", X"03", X"d0", X"04", X"d0", 
    X"05", X"d0", X"07", X"e4", X"ba", X"0a", X"04", X"bf", 
    X"00", X"01", X"04", X"fe", X"70", X"06", X"ba", X"0d", 
    X"39", X"bf", X"00", X"36", X"e5", X"25", X"45", X"26", 
    X"70", X"30", X"f5", X"71", X"75", X"72", X"10", X"f5", 
    X"73", X"90", X"00", X"15", X"75", X"f0", X"40", X"12", 
    X"0b", X"02", X"75", X"71", X"00", X"75", X"72", X"04", 
    X"75", X"73", X"00", X"90", X"00", X"27", X"75", X"f0", 
    X"40", X"12", X"0b", X"02", X"7b", X"15", X"7c", X"00", 
    X"7d", X"40", X"e4", X"f5", X"25", X"f5", X"26", X"02", 
    X"01", X"30", X"ee", X"70", X"0b", X"ba", X"0d", X"05", 
    X"bf", X"00", X"02", X"80", X"03", X"02", X"05", X"41", 
    X"c3", X"74", X"01", X"95", X"25", X"74", X"80", X"85", 
    X"26", X"f0", X"63", X"f0", X"80", X"95", X"f0", X"40", 
    X"03", X"02", X"05", X"41", X"8b", X"82", X"8c", X"83", 
    X"8d", X"f0", X"e4", X"12", X"0b", X"21", X"f5", X"33", 
    X"f5", X"34", X"f5", X"35", X"f5", X"36", X"c3", X"e5", 
    X"33", X"94", X"04", X"e5", X"34", X"64", X"80", X"94", 
    X"80", X"50", X"5d", X"e5", X"35", X"24", X"27", X"f5", 
    X"37", X"e5", X"33", X"45", X"34", X"70", X"04", X"7e", 
    X"15", X"80", X"02", X"7e", X"00", X"8e", X"38", X"75", 
    X"39", X"00", X"75", X"3a", X"40", X"75", X"3f", X"95", 
    X"75", X"40", X"15", X"75", X"41", X"80", X"85", X"38", 
    X"82", X"85", X"39", X"83", X"85", X"3a", X"f0", X"12", 
    X"0a", X"14", X"85", X"82", X"38", X"85", X"83", X"39", 
    X"85", X"f0", X"3a", X"a8", X"37", X"a6", X"38", X"08", 
    X"a6", X"39", X"08", X"a6", X"3a", X"e5", X"38", X"45", 
    X"39", X"60", X"15", X"74", X"03", X"25", X"35", X"f5", 
    X"35", X"e4", X"35", X"36", X"f5", X"36", X"05", X"33", 
    X"e4", X"b5", X"33", X"9a", X"05", X"34", X"80", X"96", 
    X"85", X"27", X"38", X"85", X"28", X"39", X"85", X"29", 
    X"3a", X"e5", X"38", X"45", X"39", X"70", X"03", X"02", 
    X"05", X"0f", X"c0", X"38", X"c0", X"39", X"c0", X"3a", 
    X"74", X"97", X"c0", X"e0", X"74", X"15", X"c0", X"e0", 
    X"74", X"80", X"c0", X"e0", X"12", X"0c", X"13", X"e5", 
    X"81", X"24", X"fa", X"f5", X"81", X"c0", X"2a", X"c0", 
    X"2b", X"c0", X"2c", X"74", X"a7", X"c0", X"e0", X"74", 
    X"15", X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", 
    X"0c", X"13", X"e5", X"81", X"24", X"fa", X"f5", X"81", 
    X"75", X"71", X"b7", X"75", X"72", X"15", X"75", X"73", 
    X"80", X"85", X"27", X"82", X"85", X"28", X"83", X"85", 
    X"29", X"f0", X"12", X"0b", X"92", X"e5", X"82", X"85", 
    X"83", X"f0", X"45", X"f0", X"70", X"58", X"85", X"2a", 
    X"38", X"85", X"2b", X"39", X"85", X"2c", X"3a", X"e5", 
    X"38", X"45", X"39", X"60", X"1e", X"85", X"38", X"82", 
    X"85", X"39", X"83", X"85", X"3a", X"f0", X"12", X"07", 
    X"94", X"85", X"82", X"38", X"85", X"83", X"39", X"ae", 
    X"38", X"53", X"06", X"0f", X"e5", X"80", X"54", X"f0", 
    X"4e", X"f5", X"80", X"85", X"80", X"38", X"75", X"39", 
    X"00", X"74", X"0f", X"55", X"38", X"f5", X"38", X"75", 
    X"39", X"00", X"c0", X"38", X"c0", X"39", X"74", X"bb", 
    X"c0", X"e0", X"74", X"15", X"c0", X"e0", X"74", X"80", 
    X"c0", X"e0", X"12", X"0c", X"13", X"e5", X"81", X"24", 
    X"fb", X"f5", X"81", X"02", X"05", X"0f", X"75", X"71", 
    X"c7", X"75", X"72", X"15", X"75", X"73", X"80", X"85", 
    X"27", X"82", X"85", X"28", X"83", X"85", X"29", X"f0", 
    X"12", X"0b", X"92", X"e5", X"82", X"85", X"83", X"f0", 
    X"45", X"f0", X"70", X"2a", X"85", X"a0", X"38", X"f5", 
    X"39", X"74", X"03", X"55", X"38", X"f5", X"38", X"75", 
    X"39", X"00", X"c0", X"38", X"c0", X"39", X"74", X"ca", 
    X"c0", X"e0", X"74", X"15", X"c0", X"e0", X"74", X"80", 
    X"c0", X"e0", X"12", X"0c", X"13", X"e5", X"81", X"24", 
    X"fb", X"f5", X"81", X"02", X"05", X"0f", X"75", X"71", 
    X"d5", X"75", X"72", X"15", X"75", X"73", X"80", X"85", 
    X"27", X"82", X"85", X"28", X"83", X"85", X"29", X"f0", 
    X"12", X"0b", X"92", X"e5", X"82", X"85", X"83", X"f0", 
    X"45", X"f0", X"70", X"21", X"85", X"08", X"38", X"f5", 
    X"39", X"c0", X"38", X"c0", X"39", X"74", X"dd", X"c0", 
    X"e0", X"74", X"15", X"c0", X"e0", X"74", X"80", X"c0", 
    X"e0", X"12", X"0c", X"13", X"e5", X"81", X"24", X"fb", 
    X"f5", X"81", X"02", X"05", X"0f", X"75", X"71", X"ed", 
    X"75", X"72", X"15", X"75", X"73", X"80", X"85", X"27", 
    X"82", X"85", X"28", X"83", X"85", X"29", X"f0", X"12", 
    X"0b", X"92", X"e5", X"82", X"85", X"83", X"f0", X"45", 
    X"f0", X"70", X"46", X"85", X"2a", X"38", X"85", X"2b", 
    X"39", X"85", X"2c", X"3a", X"e5", X"38", X"45", X"39", 
    X"60", X"15", X"85", X"38", X"82", X"85", X"39", X"83", 
    X"85", X"3a", X"f0", X"12", X"07", X"94", X"85", X"82", 
    X"38", X"85", X"83", X"39", X"85", X"38", X"80", X"85", 
    X"80", X"38", X"75", X"39", X"00", X"c0", X"38", X"c0", 
    X"39", X"74", X"f0", X"c0", X"e0", X"74", X"15", X"c0", 
    X"e0", X"74", X"80", X"c0", X"e0", X"12", X"0c", X"13", 
    X"e5", X"81", X"24", X"fb", X"f5", X"81", X"02", X"05", 
    X"0f", X"75", X"71", X"fb", X"75", X"72", X"15", X"75", 
    X"73", X"80", X"85", X"27", X"82", X"85", X"28", X"83", 
    X"85", X"29", X"f0", X"12", X"0b", X"92", X"e5", X"82", 
    X"85", X"83", X"f0", X"45", X"f0", X"70", X"46", X"85", 
    X"2a", X"38", X"85", X"2b", X"39", X"85", X"2c", X"3a", 
    X"e5", X"38", X"45", X"39", X"60", X"15", X"85", X"38", 
    X"82", X"85", X"39", X"83", X"85", X"3a", X"f0", X"12", 
    X"07", X"94", X"85", X"82", X"38", X"85", X"83", X"39", 
    X"85", X"38", X"90", X"85", X"90", X"38", X"75", X"39", 
    X"00", X"c0", X"38", X"c0", X"39", X"74", X"fe", X"c0", 
    X"e0", X"74", X"15", X"c0", X"e0", X"74", X"80", X"c0", 
    X"e0", X"12", X"0c", X"13", X"e5", X"81", X"24", X"fb", 
    X"f5", X"81", X"02", X"05", X"0f", X"75", X"71", X"09", 
    X"75", X"72", X"16", X"75", X"73", X"80", X"85", X"27", 
    X"82", X"85", X"28", X"83", X"85", X"29", X"f0", X"12", 
    X"0b", X"92", X"e5", X"82", X"85", X"83", X"f0", X"45", 
    X"f0", X"70", X"5c", X"85", X"2a", X"82", X"85", X"2b", 
    X"83", X"85", X"2c", X"f0", X"12", X"08", X"0f", X"85", 
    X"82", X"38", X"85", X"83", X"39", X"74", X"01", X"b5", 
    X"38", X"06", X"14", X"b5", X"39", X"02", X"80", X"02", 
    X"80", X"05", X"75", X"14", X"01", X"80", X"17", X"85", 
    X"2a", X"82", X"85", X"2b", X"83", X"85", X"2c", X"f0", 
    X"12", X"08", X"0f", X"e5", X"82", X"85", X"83", X"f0", 
    X"45", X"f0", X"70", X"02", X"f5", X"14", X"85", X"14", 
    X"38", X"75", X"39", X"00", X"c0", X"38", X"c0", X"39", 
    X"74", X"0f", X"c0", X"e0", X"74", X"16", X"c0", X"e0", 
    X"74", X"80", X"c0", X"e0", X"12", X"0c", X"13", X"e5", 
    X"81", X"24", X"fb", X"f5", X"81", X"80", X"38", X"85", 
    X"27", X"82", X"85", X"28", X"83", X"85", X"29", X"f0", 
    X"12", X"14", X"d9", X"60", X"2a", X"74", X"1e", X"c0", 
    X"e0", X"74", X"15", X"c0", X"e0", X"74", X"80", X"c0", 
    X"e0", X"12", X"0c", X"13", X"15", X"81", X"15", X"81", 
    X"15", X"81", X"74", X"4a", X"c0", X"e0", X"74", X"15", 
    X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", X"0c", 
    X"13", X"15", X"81", X"15", X"81", X"15", X"81", X"75", 
    X"71", X"00", X"75", X"72", X"10", X"75", X"73", X"00", 
    X"90", X"00", X"15", X"75", X"f0", X"40", X"12", X"0b", 
    X"02", X"75", X"71", X"00", X"75", X"72", X"04", X"75", 
    X"73", X"00", X"90", X"00", X"27", X"75", X"f0", X"40", 
    X"12", X"0b", X"02", X"7b", X"15", X"7c", X"00", X"7d", 
    X"40", X"e4", X"f5", X"25", X"f5", X"26", X"02", X"01", 
    X"30", X"ba", X"08", X"56", X"bf", X"00", X"53", X"c0", 
    X"05", X"c0", X"04", X"c0", X"03", X"74", X"1d", X"c0", 
    X"e0", X"74", X"16", X"c0", X"e0", X"74", X"80", X"c0", 
    X"e0", X"12", X"0c", X"13", X"15", X"81", X"15", X"81", 
    X"15", X"81", X"d0", X"03", X"d0", X"04", X"d0", X"05", 
    X"74", X"15", X"c0", X"e0", X"74", X"00", X"c0", X"e0", 
    X"74", X"40", X"c0", X"e0", X"8b", X"82", X"8c", X"83", 
    X"8d", X"f0", X"12", X"00", X"11", X"15", X"81", X"15", 
    X"81", X"15", X"81", X"70", X"03", X"02", X"01", X"30", 
    X"1b", X"bb", X"ff", X"01", X"1c", X"8b", X"82", X"8c", 
    X"83", X"8d", X"f0", X"e4", X"12", X"0b", X"21", X"02", 
    X"01", X"30", X"8b", X"82", X"8c", X"83", X"8d", X"f0", 
    X"ea", X"12", X"0b", X"21", X"a3", X"ab", X"82", X"ac", 
    X"83", X"05", X"25", X"e4", X"b5", X"25", X"02", X"05", 
    X"26", X"02", X"01", X"30", X"74", X"01", X"b5", X"14", 
    X"02", X"80", X"03", X"02", X"07", X"8a", X"74", X"f6", 
    X"25", X"08", X"40", X"3f", X"e5", X"80", X"54", X"3f", 
    X"44", X"40", X"f5", X"80", X"85", X"09", X"90", X"c0", 
    X"05", X"c0", X"04", X"c0", X"03", X"12", X"08", X"8e", 
    X"e5", X"80", X"54", X"3f", X"44", X"c0", X"f5", X"80", 
    X"e5", X"80", X"54", X"3f", X"44", X"80", X"f5", X"80", 
    X"e5", X"08", X"24", X"09", X"f9", X"87", X"90", X"12", 
    X"08", X"8e", X"d0", X"03", X"d0", X"04", X"d0", X"05", 
    X"e5", X"80", X"54", X"3f", X"44", X"c0", X"f5", X"80", 
    X"02", X"01", X"30", X"74", X"f6", X"25", X"08", X"50", 
    X"47", X"74", X"ec", X"25", X"08", X"40", X"41", X"e5", 
    X"80", X"54", X"3f", X"44", X"40", X"f5", X"80", X"85", 
    X"0a", X"90", X"c0", X"05", X"c0", X"04", X"c0", X"03", 
    X"12", X"08", X"8e", X"e5", X"80", X"54", X"3f", X"44", 
    X"c0", X"f5", X"80", X"e5", X"80", X"54", X"3f", X"44", 
    X"80", X"f5", X"80", X"e5", X"08", X"24", X"f6", X"24", 
    X"09", X"f9", X"87", X"90", X"12", X"08", X"8e", X"d0", 
    X"03", X"d0", X"04", X"d0", X"05", X"e5", X"80", X"54", 
    X"3f", X"44", X"c0", X"f5", X"80", X"02", X"01", X"30", 
    X"74", X"ec", X"25", X"08", X"50", X"47", X"74", X"e2", 
    X"25", X"08", X"40", X"41", X"e5", X"80", X"54", X"3f", 
    X"44", X"40", X"f5", X"80", X"85", X"0b", X"90", X"c0", 
    X"05", X"c0", X"04", X"c0", X"03", X"12", X"08", X"8e", 
    X"e5", X"80", X"54", X"3f", X"44", X"c0", X"f5", X"80", 
    X"e5", X"80", X"54", X"3f", X"44", X"80", X"f5", X"80", 
    X"e5", X"08", X"24", X"ec", X"24", X"09", X"f9", X"87", 
    X"90", X"12", X"08", X"8e", X"d0", X"03", X"d0", X"04", 
    X"d0", X"05", X"e5", X"80", X"54", X"3f", X"44", X"c0", 
    X"f5", X"80", X"02", X"01", X"30", X"74", X"e2", X"25", 
    X"08", X"50", X"47", X"74", X"d8", X"25", X"08", X"40", 
    X"41", X"e5", X"80", X"54", X"3f", X"44", X"40", X"f5", 
    X"80", X"85", X"0c", X"90", X"c0", X"05", X"c0", X"04", 
    X"c0", X"03", X"12", X"08", X"8e", X"e5", X"80", X"54", 
    X"3f", X"44", X"c0", X"f5", X"80", X"e5", X"80", X"54", 
    X"3f", X"44", X"80", X"f5", X"80", X"e5", X"08", X"24", 
    X"e2", X"24", X"09", X"f9", X"87", X"90", X"12", X"08", 
    X"8e", X"d0", X"03", X"d0", X"04", X"d0", X"05", X"e5", 
    X"80", X"54", X"3f", X"44", X"c0", X"f5", X"80", X"02", 
    X"01", X"30", X"74", X"d8", X"25", X"08", X"50", X"47", 
    X"74", X"ce", X"25", X"08", X"40", X"41", X"e5", X"80", 
    X"54", X"3f", X"44", X"40", X"f5", X"80", X"85", X"0d", 
    X"90", X"c0", X"05", X"c0", X"04", X"c0", X"03", X"12", 
    X"08", X"8e", X"e5", X"80", X"54", X"3f", X"44", X"c0", 
    X"f5", X"80", X"e5", X"80", X"54", X"3f", X"44", X"80", 
    X"f5", X"80", X"e5", X"08", X"24", X"d8", X"24", X"09", 
    X"f9", X"87", X"90", X"12", X"08", X"8e", X"d0", X"03", 
    X"d0", X"04", X"d0", X"05", X"e5", X"80", X"54", X"3f", 
    X"44", X"c0", X"f5", X"80", X"02", X"01", X"30", X"74", 
    X"ce", X"25", X"08", X"40", X"03", X"02", X"01", X"30", 
    X"74", X"c4", X"25", X"08", X"50", X"03", X"02", X"01", 
    X"30", X"e5", X"80", X"54", X"3f", X"44", X"40", X"f5", 
    X"80", X"85", X"0e", X"90", X"c0", X"05", X"c0", X"04", 
    X"c0", X"03", X"12", X"08", X"8e", X"e5", X"80", X"54", 
    X"3f", X"44", X"c0", X"f5", X"80", X"e5", X"80", X"54", 
    X"3f", X"44", X"80", X"f5", X"80", X"e5", X"08", X"24", 
    X"ce", X"24", X"09", X"f9", X"87", X"90", X"12", X"08", 
    X"8e", X"d0", X"03", X"d0", X"04", X"d0", X"05", X"e5", 
    X"80", X"54", X"3f", X"44", X"c0", X"f5", X"80", X"02", 
    X"01", X"30", X"53", X"80", X"3f", X"75", X"90", X"00", 
    X"02", X"01", X"30", X"22", X"ad", X"82", X"ae", X"83", 
    X"af", X"f0", X"e4", X"f5", X"71", X"f5", X"72", X"ed", 
    X"4e", X"60", X"65", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"12", X"14", X"d9", X"fa", X"60", X"59", X"ea", 
    X"24", X"c6", X"40", X"27", X"8a", X"00", X"79", X"00", 
    X"e8", X"24", X"d0", X"f8", X"e9", X"34", X"ff", X"f9", 
    X"ab", X"71", X"e5", X"72", X"c4", X"54", X"f0", X"cb", 
    X"c4", X"cb", X"6b", X"cb", X"54", X"f0", X"cb", X"6b", 
    X"fc", X"eb", X"28", X"f5", X"71", X"ec", X"39", X"f5", 
    X"72", X"80", X"26", X"53", X"02", X"5f", X"7c", X"00", 
    X"74", X"c9", X"2a", X"fa", X"74", X"ff", X"3c", X"fc", 
    X"ab", X"71", X"e5", X"72", X"c4", X"54", X"f0", X"cb", 
    X"c4", X"cb", X"6b", X"cb", X"54", X"f0", X"cb", X"6b", 
    X"f9", X"eb", X"2a", X"f5", X"71", X"e9", X"3c", X"f5", 
    X"72", X"0d", X"bd", X"00", X"9a", X"0e", X"80", X"97", 
    X"85", X"71", X"82", X"85", X"72", X"83", X"22", X"ad", 
    X"82", X"ae", X"83", X"af", X"f0", X"e4", X"f5", X"71", 
    X"f5", X"72", X"f5", X"73", X"f5", X"74", X"ed", X"4e", 
    X"60", X"52", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"14", X"d9", X"f8", X"60", X"46", X"b8", X"2d", 
    X"08", X"75", X"73", X"01", X"75", X"74", X"00", X"80", 
    X"34", X"7a", X"00", X"e8", X"24", X"d0", X"f8", X"ea", 
    X"34", X"ff", X"fa", X"a9", X"71", X"e5", X"72", X"c4", 
    X"03", X"54", X"f8", X"c9", X"c4", X"03", X"c9", X"69", 
    X"c9", X"54", X"f8", X"c9", X"69", X"fc", X"e9", X"28", 
    X"f8", X"ec", X"3a", X"fa", X"e5", X"71", X"25", X"71", 
    X"fb", X"e5", X"72", X"33", X"fc", X"eb", X"28", X"f5", 
    X"71", X"ec", X"3a", X"f5", X"72", X"0d", X"bd", X"00", 
    X"ad", X"0e", X"80", X"aa", X"e5", X"73", X"45", X"74", 
    X"60", X"0b", X"c3", X"e4", X"95", X"71", X"fe", X"e4", 
    X"95", X"72", X"ff", X"80", X"04", X"ae", X"71", X"af", 
    X"72", X"8e", X"82", X"8f", X"83", X"22", X"7e", X"88", 
    X"7f", X"13", X"ee", X"24", X"ff", X"fc", X"ef", X"34", 
    X"ff", X"fd", X"8c", X"06", X"8d", X"07", X"ec", X"4d", 
    X"70", X"f0", X"22", X"75", X"08", X"00", X"90", X"c3", 
    X"50", X"12", X"09", X"29", X"75", X"82", X"01", X"12", 
    X"09", X"76", X"75", X"82", X"01", X"12", X"09", X"20", 
    X"75", X"82", X"01", X"12", X"09", X"46", X"22", X"12", 
    X"09", X"4f", X"ae", X"82", X"af", X"83", X"7d", X"00", 
    X"7c", X"00", X"75", X"71", X"32", X"e4", X"f5", X"72", 
    X"f5", X"73", X"f5", X"74", X"8e", X"82", X"8f", X"83", 
    X"8d", X"f0", X"ec", X"12", X"09", X"af", X"ac", X"82", 
    X"ad", X"83", X"ae", X"f0", X"ff", X"85", X"08", X"71", 
    X"75", X"72", X"00", X"90", X"03", X"e8", X"c0", X"07", 
    X"c0", X"06", X"c0", X"05", X"c0", X"04", X"12", X"0b", 
    X"75", X"aa", X"82", X"ab", X"83", X"d0", X"04", X"d0", 
    X"05", X"d0", X"06", X"d0", X"07", X"8a", X"00", X"eb", 
    X"f9", X"33", X"95", X"e0", X"fa", X"fb", X"e8", X"2c", 
    X"fc", X"e9", X"3d", X"fd", X"ea", X"3e", X"fe", X"eb", 
    X"3f", X"8c", X"82", X"8d", X"83", X"8e", X"f0", X"22", 
    X"e5", X"82", X"54", X"01", X"24", X"ff", X"92", X"af", 
    X"22", X"ae", X"82", X"af", X"83", X"8e", X"04", X"8f", 
    X"05", X"bc", X"ff", X"05", X"bd", X"ff", X"02", X"80", 
    X"08", X"8f", X"8f", X"8e", X"8e", X"d2", X"8c", X"80", 
    X"02", X"c2", X"8c", X"d2", X"88", X"22", X"e5", X"82", 
    X"54", X"01", X"24", X"ff", X"92", X"8d", X"22", X"85", 
    X"8d", X"71", X"85", X"8c", X"72", X"85", X"8c", X"73", 
    X"e5", X"73", X"b5", X"72", X"02", X"80", X"06", X"85", 
    X"8d", X"71", X"85", X"8c", X"72", X"af", X"71", X"7e", 
    X"00", X"ac", X"72", X"7d", X"00", X"ec", X"4e", X"f5", 
    X"82", X"ed", X"4f", X"f5", X"83", X"22", X"e5", X"82", 
    X"54", X"01", X"24", X"ff", X"92", X"a9", X"22", X"c0", 
    X"e0", X"c0", X"d0", X"d2", X"88", X"05", X"3b", X"74", 
    X"3b", X"b5", X"08", X"05", X"75", X"08", X"00", X"80", 
    X"05", X"e5", X"08", X"04", X"f5", X"08", X"d0", X"d0", 
    X"d0", X"e0", X"32", X"ae", X"82", X"30", X"9c", X"fd", 
    X"8e", X"99", X"22", X"30", X"9d", X"fd", X"ae", X"99", 
    X"7f", X"00", X"8e", X"82", X"8f", X"83", X"22", X"fb", 
    X"7a", X"20", X"e4", X"fc", X"fd", X"fe", X"ff", X"e5", 
    X"82", X"25", X"82", X"f5", X"82", X"e5", X"83", X"33", 
    X"f5", X"83", X"e5", X"f0", X"33", X"f5", X"f0", X"eb", 
    X"33", X"fb", X"40", X"17", X"da", X"e9", X"80", X"42", 
    X"e5", X"82", X"25", X"82", X"f5", X"82", X"e5", X"83", 
    X"33", X"f5", X"83", X"e5", X"f0", X"33", X"f5", X"f0", 
    X"eb", X"33", X"fb", X"ec", X"33", X"fc", X"ed", X"33", 
    X"fd", X"ee", X"33", X"fe", X"ef", X"33", X"ff", X"ec", 
    X"95", X"71", X"ed", X"95", X"72", X"ee", X"95", X"73", 
    X"ef", X"95", X"74", X"40", X"13", X"ec", X"95", X"71", 
    X"fc", X"ed", X"95", X"72", X"fd", X"ee", X"95", X"73", 
    X"fe", X"ef", X"95", X"74", X"ff", X"43", X"82", X"01", 
    X"da", X"be", X"eb", X"22", X"ad", X"82", X"ae", X"83", 
    X"af", X"f0", X"ed", X"4e", X"60", X"06", X"8d", X"3c", 
    X"8e", X"3d", X"8f", X"3e", X"e5", X"3c", X"45", X"3d", 
    X"70", X"06", X"90", X"00", X"00", X"f5", X"f0", X"22", 
    X"ad", X"3c", X"ae", X"3d", X"af", X"3e", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"12", X"14", X"d9", X"60", 
    X"31", X"ad", X"3c", X"ae", X"3d", X"af", X"3e", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"14", X"d9", 
    X"f5", X"71", X"85", X"3f", X"82", X"85", X"40", X"83", 
    X"85", X"41", X"f0", X"12", X"0b", X"3c", X"ad", X"82", 
    X"ae", X"83", X"af", X"f0", X"ed", X"4e", X"60", X"0a", 
    X"05", X"3c", X"e4", X"b5", X"3c", X"c2", X"05", X"3d", 
    X"80", X"be", X"ad", X"3c", X"ae", X"3d", X"af", X"3e", 
    X"aa", X"3c", X"ab", X"3d", X"ac", X"3e", X"8a", X"82", 
    X"8b", X"83", X"8c", X"f0", X"12", X"14", X"d9", X"60", 
    X"59", X"aa", X"3c", X"ab", X"3d", X"ac", X"3e", X"8a", 
    X"82", X"8b", X"83", X"8c", X"f0", X"12", X"14", X"d9", 
    X"f5", X"71", X"85", X"3f", X"82", X"85", X"40", X"83", 
    X"85", X"41", X"f0", X"c0", X"07", X"c0", X"06", X"c0", 
    X"05", X"12", X"0b", X"3c", X"aa", X"82", X"ab", X"83", 
    X"d0", X"05", X"d0", X"06", X"d0", X"07", X"ea", X"4b", 
    X"60", X"1e", X"aa", X"3c", X"ab", X"3d", X"ac", X"3e", 
    X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"e4", X"12", 
    X"0b", X"21", X"05", X"3c", X"b5", X"3c", X"02", X"05", 
    X"3d", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"22", 
    X"05", X"3c", X"e4", X"b5", X"3c", X"9a", X"05", X"3d", 
    X"80", X"96", X"e4", X"f5", X"3c", X"f5", X"3d", X"f5", 
    X"3e", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", 
    X"14", X"d9", X"60", X"07", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"22", X"90", X"00", X"00", X"75", X"f0", 
    X"00", X"22", X"ac", X"82", X"ad", X"83", X"ae", X"72", 
    X"af", X"73", X"be", X"00", X"04", X"ef", X"60", X"0c", 
    X"1f", X"0f", X"e5", X"71", X"12", X"0b", X"21", X"a3", 
    X"de", X"fa", X"df", X"f8", X"8c", X"82", X"8d", X"83", 
    X"22", X"20", X"f7", X"11", X"30", X"f6", X"13", X"88", 
    X"83", X"a8", X"82", X"20", X"f5", X"09", X"f6", X"a8", 
    X"83", X"75", X"83", X"00", X"22", X"80", X"fe", X"f2", 
    X"80", X"f5", X"f0", X"22", X"ad", X"82", X"ae", X"83", 
    X"af", X"f0", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"14", X"d9", X"fc", X"60", X"0d", X"ec", X"b5", 
    X"71", X"02", X"80", X"07", X"0d", X"bd", X"00", X"ea", 
    X"0e", X"80", X"e7", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"12", X"14", X"d9", X"b5", X"71", X"07", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"22", X"90", X"00", 
    X"00", X"75", X"f0", X"00", X"22", X"e5", X"82", X"85", 
    X"71", X"f0", X"a4", X"c5", X"82", X"c0", X"f0", X"85", 
    X"72", X"f0", X"a4", X"d0", X"f0", X"25", X"f0", X"c5", 
    X"83", X"85", X"71", X"f0", X"a4", X"25", X"83", X"f5", 
    X"83", X"22", X"ad", X"82", X"ae", X"83", X"af", X"f0", 
    X"aa", X"71", X"ab", X"72", X"ac", X"73", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"12", X"14", X"d9", X"f8", 
    X"79", X"00", X"8a", X"82", X"8b", X"83", X"8c", X"f0", 
    X"12", X"14", X"d9", X"f5", X"74", X"c0", X"02", X"c0", 
    X"03", X"c0", X"04", X"ab", X"74", X"7c", X"00", X"e8", 
    X"c3", X"9b", X"f8", X"e9", X"9c", X"f9", X"88", X"75", 
    X"89", X"76", X"d0", X"04", X"d0", X"03", X"d0", X"02", 
    X"e8", X"49", X"70", X"10", X"e5", X"74", X"60", X"0c", 
    X"0d", X"bd", X"00", X"01", X"0e", X"0a", X"ba", X"00", 
    X"bd", X"0b", X"80", X"ba", X"85", X"75", X"82", X"85", 
    X"76", X"83", X"22", X"c0", X"70", X"85", X"81", X"70", 
    X"7e", X"00", X"8e", X"83", X"12", X"09", X"9b", X"d0", 
    X"70", X"22", X"85", X"82", X"53", X"85", X"83", X"54", 
    X"85", X"f0", X"55", X"e4", X"f5", X"50", X"f5", X"51", 
    X"f5", X"52", X"85", X"42", X"56", X"90", X"0b", X"eb", 
    X"02", X"0c", X"d9", X"c0", X"70", X"e5", X"81", X"f5", 
    X"70", X"24", X"fb", X"ff", X"8f", X"56", X"e4", X"f5", 
    X"50", X"f5", X"51", X"f5", X"52", X"e5", X"70", X"24", 
    X"fb", X"f8", X"86", X"53", X"08", X"86", X"54", X"08", 
    X"86", X"55", X"90", X"0b", X"eb", X"12", X"0c", X"d9", 
    X"d0", X"70", X"22", X"af", X"82", X"c0", X"46", X"c0", 
    X"47", X"c0", X"48", X"12", X"0c", X"48", X"80", X"07", 
    X"c0", X"44", X"c0", X"45", X"8f", X"82", X"22", X"15", 
    X"81", X"15", X"81", X"15", X"81", X"05", X"4e", X"e4", 
    X"b5", X"4e", X"02", X"05", X"4f", X"22", X"af", X"82", 
    X"74", X"30", X"2f", X"ff", X"24", X"c6", X"50", X"0b", 
    X"74", X"07", X"2f", X"ff", X"e5", X"43", X"60", X"03", 
    X"43", X"07", X"20", X"8f", X"82", X"02", X"0c", X"3b", 
    X"e5", X"82", X"ff", X"c4", X"54", X"0f", X"f5", X"82", 
    X"c0", X"07", X"12", X"0c", X"5e", X"d0", X"07", X"74", 
    X"0f", X"5f", X"f5", X"82", X"02", X"0c", X"5e", X"85", 
    X"82", X"71", X"ab", X"49", X"ac", X"4a", X"ad", X"4b", 
    X"ae", X"4c", X"aa", X"4d", X"75", X"73", X"20", X"8a", 
    X"07", X"ef", X"2f", X"f5", X"72", X"ee", X"23", X"54", 
    X"01", X"45", X"72", X"fa", X"eb", X"2b", X"fb", X"ec", 
    X"33", X"fc", X"ed", X"33", X"fd", X"ee", X"33", X"fe", 
    X"c3", X"ea", X"95", X"71", X"40", X"08", X"ea", X"c3", 
    X"95", X"71", X"fa", X"43", X"03", X"01", X"e5", X"73", 
    X"14", X"ff", X"8f", X"73", X"70", X"d1", X"8b", X"49", 
    X"8c", X"4a", X"8d", X"4b", X"8e", X"4c", X"8a", X"4d", 
    X"22", X"85", X"82", X"44", X"85", X"83", X"45", X"85", 
    X"50", X"46", X"85", X"51", X"47", X"85", X"52", X"48", 
    X"e4", X"f5", X"4e", X"f5", X"4f", X"ad", X"53", X"ae", 
    X"54", X"af", X"55", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"12", X"14", X"d9", X"fc", X"74", X"01", X"2d", 
    X"f5", X"53", X"e4", X"3e", X"f5", X"54", X"8f", X"55", 
    X"ec", X"ff", X"70", X"03", X"02", X"14", X"ba", X"bf", 
    X"25", X"02", X"80", X"03", X"02", X"14", X"b2", X"7e", 
    X"00", X"7d", X"00", X"8e", X"57", X"8e", X"58", X"7a", 
    X"00", X"7b", X"00", X"8e", X"59", X"7c", X"00", X"8e", 
    X"5a", X"e4", X"f5", X"62", X"f5", X"63", X"75", X"5b", 
    X"ff", X"75", X"5c", X"ff", X"85", X"53", X"64", X"85", 
    X"54", X"65", X"85", X"55", X"66", X"85", X"64", X"82", 
    X"85", X"65", X"83", X"85", X"66", X"f0", X"12", X"14", 
    X"d9", X"f5", X"67", X"a3", X"85", X"82", X"64", X"85", 
    X"83", X"65", X"85", X"64", X"53", X"85", X"65", X"54", 
    X"85", X"66", X"55", X"74", X"25", X"b5", X"67", X"08", 
    X"85", X"67", X"82", X"12", X"0c", X"3b", X"80", X"85", 
    X"74", X"d0", X"25", X"67", X"40", X"03", X"02", X"0e", 
    X"1b", X"e5", X"67", X"24", X"c6", X"50", X"03", X"02", 
    X"0e", X"1b", X"74", X"ff", X"b5", X"5b", X"55", X"b5", 
    X"5c", X"52", X"85", X"62", X"71", X"85", X"63", X"72", 
    X"90", X"00", X"0a", X"c0", X"06", X"c0", X"05", X"c0", 
    X"04", X"c0", X"03", X"c0", X"02", X"12", X"0b", X"75", 
    X"85", X"82", X"68", X"85", X"83", X"69", X"d0", X"02", 
    X"d0", X"03", X"d0", X"04", X"d0", X"05", X"d0", X"06", 
    X"85", X"67", X"6a", X"75", X"6b", X"00", X"e5", X"6a", 
    X"25", X"68", X"f5", X"6a", X"e5", X"6b", X"35", X"69", 
    X"f5", X"6b", X"e5", X"6a", X"24", X"d0", X"f5", X"62", 
    X"e5", X"6b", X"34", X"ff", X"f5", X"63", X"e5", X"62", 
    X"45", X"63", X"60", X"03", X"02", X"0d", X"3d", X"7d", 
    X"01", X"02", X"0d", X"3d", X"85", X"5b", X"71", X"85", 
    X"5c", X"72", X"90", X"00", X"0a", X"c0", X"06", X"c0", 
    X"05", X"c0", X"04", X"c0", X"03", X"c0", X"02", X"12", 
    X"0b", X"75", X"85", X"82", X"6a", X"85", X"83", X"6b", 
    X"d0", X"02", X"d0", X"03", X"d0", X"04", X"d0", X"05", 
    X"d0", X"06", X"85", X"67", X"68", X"75", X"69", X"00", 
    X"e5", X"68", X"25", X"6a", X"f5", X"6a", X"e5", X"69", 
    X"35", X"6b", X"f5", X"6b", X"e5", X"6a", X"24", X"d0", 
    X"f5", X"5b", X"e5", X"6b", X"34", X"ff", X"f5", X"5c", 
    X"02", X"0d", X"3d", X"74", X"2e", X"b5", X"67", X"15", 
    X"74", X"ff", X"b5", X"5b", X"05", X"b5", X"5c", X"02", 
    X"80", X"03", X"02", X"0d", X"3d", X"e4", X"f5", X"5b", 
    X"f5", X"5c", X"02", X"0d", X"3d", X"74", X"9f", X"25", 
    X"67", X"50", X"0e", X"e5", X"67", X"24", X"85", X"40", 
    X"08", X"53", X"67", X"df", X"75", X"43", X"01", X"80", 
    X"03", X"75", X"43", X"00", X"74", X"20", X"b5", X"67", 
    X"03", X"02", X"0e", X"e7", X"74", X"2b", X"b5", X"67", 
    X"03", X"02", X"0e", X"e1", X"74", X"2d", X"b5", X"67", 
    X"02", X"80", X"79", X"74", X"42", X"b5", X"67", X"03", 
    X"02", X"0e", X"ed", X"74", X"43", X"b5", X"67", X"03", 
    X"02", X"0e", X"f8", X"74", X"44", X"b5", X"67", X"03", 
    X"02", X"11", X"45", X"74", X"46", X"b5", X"67", X"03", 
    X"02", X"11", X"5b", X"74", X"48", X"b5", X"67", X"03", 
    X"02", X"0d", X"3d", X"74", X"49", X"b5", X"67", X"03", 
    X"02", X"11", X"45", X"74", X"4a", X"b5", X"67", X"03", 
    X"02", X"0d", X"3d", X"74", X"4c", X"b5", X"67", X"02", 
    X"80", X"50", X"74", X"4f", X"b5", X"67", X"03", X"02", 
    X"11", X"4c", X"74", X"50", X"b5", X"67", X"03", X"02", 
    X"10", X"90", X"74", X"53", X"b5", X"67", X"02", X"80", 
    X"76", X"74", X"54", X"b5", X"67", X"03", X"02", X"0d", 
    X"3d", X"74", X"55", X"b5", X"67", X"03", X"02", X"11", 
    X"51", X"74", X"58", X"b5", X"67", X"03", X"02", X"11", 
    X"56", X"74", X"5a", X"b5", X"67", X"03", X"02", X"0d", 
    X"3d", X"02", X"11", X"5f", X"7e", X"01", X"02", X"0d", 
    X"3d", X"75", X"57", X"01", X"02", X"0d", X"3d", X"75", 
    X"58", X"01", X"02", X"0d", X"3d", X"7b", X"01", X"02", 
    X"0d", X"3d", X"75", X"59", X"01", X"02", X"0d", X"3d", 
    X"eb", X"60", X"0a", X"e5", X"56", X"14", X"f9", X"89", 
    X"56", X"87", X"6a", X"80", X"0d", X"e5", X"56", X"24", 
    X"fe", X"f5", X"68", X"85", X"68", X"56", X"a9", X"68", 
    X"87", X"6a", X"85", X"6a", X"82", X"c0", X"06", X"c0", 
    X"05", X"c0", X"04", X"c0", X"03", X"c0", X"02", X"12", 
    X"0c", X"3b", X"d0", X"02", X"d0", X"03", X"d0", X"04", 
    X"d0", X"05", X"d0", X"06", X"02", X"11", X"81", X"e5", 
    X"56", X"24", X"fd", X"f5", X"6a", X"85", X"6a", X"56", 
    X"a9", X"6a", X"87", X"64", X"09", X"87", X"65", X"09", 
    X"87", X"66", X"19", X"19", X"85", X"64", X"49", X"85", 
    X"65", X"4a", X"85", X"66", X"4b", X"85", X"64", X"82", 
    X"85", X"65", X"83", X"85", X"66", X"f0", X"c0", X"06", 
    X"c0", X"05", X"c0", X"04", X"c0", X"03", X"c0", X"02", 
    X"12", X"14", X"c1", X"85", X"82", X"6a", X"85", X"83", 
    X"6b", X"d0", X"02", X"d0", X"03", X"d0", X"04", X"d0", 
    X"05", X"d0", X"06", X"74", X"ff", X"b5", X"5b", X"09", 
    X"b5", X"5c", X"06", X"85", X"6a", X"5b", X"85", X"6b", 
    X"5c", X"ee", X"70", X"4f", X"c3", X"e5", X"6a", X"95", 
    X"62", X"e5", X"6b", X"95", X"63", X"50", X"44", X"e5", 
    X"62", X"c3", X"95", X"6a", X"f5", X"68", X"e5", X"63", 
    X"95", X"6b", X"f5", X"69", X"85", X"68", X"64", X"85", 
    X"69", X"65", X"15", X"68", X"74", X"ff", X"b5", X"68", 
    X"02", X"15", X"69", X"e5", X"64", X"45", X"65", X"60", 
    X"1c", X"75", X"82", X"20", X"c0", X"06", X"c0", X"05", 
    X"c0", X"04", X"c0", X"03", X"c0", X"02", X"12", X"0c", 
    X"3b", X"d0", X"02", X"d0", X"03", X"d0", X"04", X"d0", 
    X"05", X"d0", X"06", X"80", X"cf", X"85", X"68", X"62", 
    X"85", X"69", X"63", X"85", X"5b", X"68", X"85", X"5c", 
    X"69", X"85", X"49", X"82", X"85", X"4a", X"83", X"85", 
    X"4b", X"f0", X"12", X"14", X"d9", X"f5", X"64", X"85", 
    X"64", X"5f", X"60", X"4f", X"c3", X"e4", X"95", X"68", 
    X"74", X"80", X"85", X"69", X"f0", X"63", X"f0", X"80", 
    X"95", X"f0", X"50", X"3f", X"15", X"68", X"74", X"ff", 
    X"b5", X"68", X"02", X"15", X"69", X"85", X"5f", X"82", 
    X"c0", X"06", X"c0", X"05", X"c0", X"04", X"c0", X"03", 
    X"c0", X"02", X"12", X"0c", X"3b", X"d0", X"02", X"d0", 
    X"03", X"d0", X"04", X"d0", X"05", X"d0", X"06", X"85", 
    X"49", X"64", X"85", X"4a", X"65", X"85", X"4b", X"66", 
    X"05", X"64", X"e4", X"b5", X"64", X"02", X"05", X"65", 
    X"85", X"64", X"49", X"85", X"65", X"4a", X"85", X"66", 
    X"4b", X"80", X"9e", X"ee", X"70", X"03", X"02", X"11", 
    X"81", X"c3", X"e5", X"6a", X"95", X"62", X"e5", X"6b", 
    X"95", X"63", X"40", X"03", X"02", X"11", X"81", X"e5", 
    X"62", X"c3", X"95", X"6a", X"f5", X"6a", X"e5", X"63", 
    X"95", X"6b", X"f5", X"6b", X"85", X"6a", X"68", X"85", 
    X"6b", X"69", X"15", X"6a", X"74", X"ff", X"b5", X"6a", 
    X"02", X"15", X"6b", X"e5", X"68", X"45", X"69", X"70", 
    X"03", X"02", X"11", X"7b", X"75", X"82", X"20", X"c0", 
    X"06", X"c0", X"05", X"c0", X"04", X"c0", X"03", X"c0", 
    X"02", X"12", X"0c", X"3b", X"d0", X"02", X"d0", X"03", 
    X"d0", X"04", X"d0", X"05", X"d0", X"06", X"80", X"cc", 
    X"e5", X"56", X"24", X"fd", X"f5", X"68", X"85", X"68", 
    X"56", X"a9", X"68", X"87", X"64", X"09", X"87", X"65", 
    X"09", X"87", X"66", X"19", X"19", X"85", X"64", X"49", 
    X"85", X"65", X"4a", X"85", X"66", X"4b", X"85", X"4b", 
    X"60", X"74", X"80", X"25", X"60", X"50", X"05", X"75", 
    X"68", X"43", X"80", X"19", X"74", X"a0", X"25", X"60", 
    X"50", X"05", X"75", X"68", X"50", X"80", X"0e", X"74", 
    X"c0", X"25", X"60", X"50", X"05", X"75", X"68", X"49", 
    X"80", X"03", X"75", X"68", X"58", X"85", X"68", X"82", 
    X"c0", X"06", X"c0", X"05", X"c0", X"04", X"c0", X"03", 
    X"c0", X"02", X"12", X"0c", X"3b", X"75", X"82", X"3a", 
    X"12", X"0c", X"3b", X"75", X"82", X"30", X"12", X"0c", 
    X"3b", X"75", X"82", X"78", X"12", X"0c", X"3b", X"d0", 
    X"02", X"d0", X"03", X"d0", X"04", X"d0", X"05", X"d0", 
    X"06", X"74", X"49", X"b5", X"68", X"02", X"80", X"21", 
    X"74", X"50", X"b5", X"68", X"02", X"80", X"1a", X"85", 
    X"4a", X"82", X"c0", X"06", X"c0", X"05", X"c0", X"04", 
    X"c0", X"03", X"c0", X"02", X"12", X"0c", X"78", X"d0", 
    X"02", X"d0", X"03", X"d0", X"04", X"d0", X"05", X"d0", 
    X"06", X"85", X"49", X"82", X"c0", X"06", X"c0", X"05", 
    X"c0", X"04", X"c0", X"03", X"c0", X"02", X"12", X"0c", 
    X"78", X"d0", X"02", X"d0", X"03", X"d0", X"04", X"d0", 
    X"05", X"d0", X"06", X"80", X"3c", X"7a", X"01", X"75", 
    X"5a", X"0a", X"80", X"35", X"75", X"5a", X"08", X"80", 
    X"30", X"75", X"5a", X"0a", X"80", X"2b", X"75", X"5a", 
    X"10", X"80", X"26", X"7c", X"01", X"80", X"22", X"85", 
    X"67", X"82", X"c0", X"06", X"c0", X"05", X"c0", X"04", 
    X"c0", X"03", X"c0", X"02", X"12", X"0c", X"3b", X"d0", 
    X"02", X"d0", X"03", X"d0", X"04", X"d0", X"05", X"d0", 
    X"06", X"80", X"06", X"85", X"6a", X"62", X"85", X"6b", 
    X"63", X"ec", X"60", X"68", X"e5", X"56", X"24", X"fc", 
    X"fc", X"8c", X"56", X"8c", X"01", X"87", X"6c", X"09", 
    X"87", X"6d", X"09", X"87", X"6e", X"09", X"87", X"6f", 
    X"19", X"19", X"19", X"85", X"6c", X"49", X"85", X"6d", 
    X"4a", X"85", X"6e", X"4b", X"85", X"6f", X"4c", X"75", 
    X"49", X"2a", X"75", X"4a", X"16", X"75", X"4b", X"80", 
    X"85", X"49", X"6c", X"85", X"4a", X"6d", X"85", X"4b", 
    X"6e", X"74", X"01", X"25", X"6c", X"f5", X"64", X"e4", 
    X"35", X"6d", X"f5", X"65", X"85", X"6e", X"66", X"85", 
    X"64", X"49", X"85", X"65", X"4a", X"85", X"66", X"4b", 
    X"85", X"6c", X"82", X"85", X"6d", X"83", X"85", X"6e", 
    X"f0", X"12", X"14", X"d9", X"fc", X"8c", X"6c", X"70", 
    X"03", X"02", X"0c", X"ed", X"85", X"6c", X"82", X"12", 
    X"0c", X"3b", X"80", X"c4", X"e5", X"5a", X"70", X"03", 
    X"02", X"0c", X"ed", X"eb", X"60", X"3f", X"e5", X"56", 
    X"14", X"f9", X"89", X"56", X"87", X"04", X"8c", X"6c", 
    X"75", X"6d", X"00", X"75", X"6e", X"00", X"75", X"6f", 
    X"00", X"85", X"6c", X"49", X"85", X"6d", X"4a", X"85", 
    X"6e", X"4b", X"85", X"6f", X"4c", X"ea", X"60", X"03", 
    X"02", X"12", X"9e", X"85", X"49", X"6c", X"75", X"6d", 
    X"00", X"75", X"6e", X"00", X"75", X"6f", X"00", X"85", 
    X"6c", X"49", X"85", X"6d", X"4a", X"85", X"6e", X"4b", 
    X"85", X"6f", X"4c", X"80", X"69", X"e5", X"59", X"60", 
    X"25", X"e5", X"56", X"24", X"fc", X"fc", X"8c", X"56", 
    X"8c", X"01", X"87", X"6c", X"09", X"87", X"6d", X"09", 
    X"87", X"6e", X"09", X"87", X"6f", X"19", X"19", X"19", 
    X"85", X"6c", X"49", X"85", X"6d", X"4a", X"85", X"6e", 
    X"4b", X"85", X"6f", X"4c", X"80", X"40", X"e5", X"56", 
    X"24", X"fe", X"fc", X"8c", X"56", X"8c", X"01", X"87", 
    X"03", X"09", X"87", X"04", X"19", X"8b", X"6c", X"ec", 
    X"f5", X"6d", X"33", X"95", X"e0", X"f5", X"6e", X"f5", 
    X"6f", X"85", X"6c", X"49", X"85", X"6d", X"4a", X"85", 
    X"6e", X"4b", X"85", X"6f", X"4c", X"ea", X"70", X"16", 
    X"85", X"49", X"6c", X"85", X"4a", X"6d", X"f5", X"6e", 
    X"f5", X"6f", X"85", X"6c", X"49", X"85", X"6d", X"4a", 
    X"85", X"6e", X"4b", X"85", X"6f", X"4c", X"ea", X"60", 
    X"2a", X"e5", X"4c", X"30", X"e7", X"23", X"c3", X"e4", 
    X"95", X"49", X"f5", X"6c", X"e4", X"95", X"4a", X"f5", 
    X"6d", X"e4", X"95", X"4b", X"f5", X"6e", X"e4", X"95", 
    X"4c", X"f5", X"6f", X"85", X"6c", X"49", X"85", X"6d", 
    X"4a", X"85", X"6e", X"4b", X"85", X"6f", X"4c", X"80", 
    X"02", X"7a", X"00", X"7c", X"01", X"79", X"7c", X"e4", 
    X"f5", X"6c", X"f5", X"6d", X"75", X"4d", X"00", X"85", 
    X"5a", X"82", X"c0", X"06", X"c0", X"05", X"c0", X"04", 
    X"c0", X"02", X"c0", X"01", X"12", X"0c", X"8f", X"d0", 
    X"01", X"d0", X"02", X"d0", X"04", X"d0", X"05", X"d0", 
    X"06", X"ec", X"70", X"0d", X"e5", X"4d", X"c4", X"f5", 
    X"6a", X"e7", X"fb", X"45", X"6a", X"f7", X"19", X"80", 
    X"02", X"a7", X"4d", X"05", X"6c", X"e4", X"b5", X"6c", 
    X"02", X"05", X"6d", X"ec", X"b4", X"01", X"00", X"e4", 
    X"33", X"fc", X"e5", X"49", X"45", X"4a", X"45", X"4b", 
    X"45", X"4c", X"70", X"b8", X"89", X"61", X"85", X"6c", 
    X"5d", X"85", X"6d", X"5e", X"e5", X"62", X"45", X"63", 
    X"70", X"05", X"75", X"62", X"01", X"f5", X"63", X"ed", 
    X"70", X"43", X"ee", X"70", X"40", X"85", X"62", X"6c", 
    X"85", X"63", X"6d", X"ab", X"5d", X"0b", X"8b", X"6a", 
    X"75", X"6b", X"00", X"c3", X"e5", X"6a", X"95", X"6c", 
    X"e5", X"6b", X"95", X"6d", X"50", X"21", X"75", X"82", 
    X"20", X"c0", X"06", X"c0", X"05", X"c0", X"04", X"c0", 
    X"02", X"12", X"0c", X"3b", X"d0", X"02", X"d0", X"04", 
    X"d0", X"05", X"d0", X"06", X"15", X"6c", X"74", X"ff", 
    X"b5", X"6c", X"02", X"15", X"6d", X"80", X"cc", X"85", 
    X"6c", X"62", X"85", X"6d", X"63", X"ea", X"60", X"1d", 
    X"75", X"82", X"2d", X"c0", X"06", X"c0", X"05", X"c0", 
    X"04", X"12", X"0c", X"3b", X"d0", X"04", X"d0", X"05", 
    X"d0", X"06", X"15", X"62", X"74", X"ff", X"b5", X"62", 
    X"02", X"15", X"63", X"80", X"46", X"e5", X"5d", X"45", 
    X"5e", X"60", X"40", X"e5", X"57", X"60", X"1d", X"75", 
    X"82", X"2b", X"c0", X"06", X"c0", X"05", X"c0", X"04", 
    X"12", X"0c", X"3b", X"d0", X"04", X"d0", X"05", X"d0", 
    X"06", X"15", X"62", X"74", X"ff", X"b5", X"62", X"02", 
    X"15", X"63", X"80", X"1f", X"e5", X"58", X"60", X"1b", 
    X"75", X"82", X"20", X"c0", X"06", X"c0", X"05", X"c0", 
    X"04", X"12", X"0c", X"3b", X"d0", X"04", X"d0", X"05", 
    X"d0", X"06", X"15", X"62", X"74", X"ff", X"b5", X"62", 
    X"02", X"15", X"63", X"ee", X"70", X"3c", X"85", X"62", 
    X"6c", X"85", X"63", X"6d", X"aa", X"6c", X"ab", X"6d", 
    X"15", X"6c", X"74", X"ff", X"b5", X"6c", X"02", X"15", 
    X"6d", X"c3", X"e5", X"5d", X"9a", X"e5", X"5e", X"9b", 
    X"50", X"41", X"ed", X"60", X"06", X"7a", X"30", X"7b", 
    X"00", X"80", X"04", X"7a", X"20", X"7b", X"00", X"8a", 
    X"82", X"c0", X"06", X"c0", X"05", X"c0", X"04", X"12", 
    X"0c", X"3b", X"d0", X"04", X"d0", X"05", X"d0", X"06", 
    X"80", X"ca", X"c3", X"e5", X"5d", X"95", X"62", X"e5", 
    X"5e", X"95", X"63", X"50", X"0f", X"e5", X"62", X"c3", 
    X"95", X"5d", X"f5", X"6a", X"e5", X"63", X"95", X"5e", 
    X"f5", X"6b", X"80", X"0d", X"e4", X"f5", X"6a", X"f5", 
    X"6b", X"80", X"06", X"85", X"6c", X"6a", X"85", X"6d", 
    X"6b", X"a9", X"61", X"85", X"5d", X"6c", X"85", X"5e", 
    X"6d", X"aa", X"6c", X"ad", X"6d", X"15", X"6c", X"74", 
    X"ff", X"b5", X"6c", X"02", X"15", X"6d", X"ea", X"4d", 
    X"60", X"2e", X"ec", X"b4", X"01", X"00", X"e4", X"33", 
    X"fc", X"70", X"0a", X"09", X"e7", X"c4", X"54", X"0f", 
    X"fd", X"8d", X"4d", X"80", X"07", X"87", X"05", X"74", 
    X"0f", X"5d", X"f5", X"4d", X"85", X"4d", X"82", X"c0", 
    X"06", X"c0", X"04", X"c0", X"01", X"12", X"0c", X"5e", 
    X"d0", X"01", X"d0", X"04", X"d0", X"06", X"80", X"c1", 
    X"ee", X"70", X"03", X"02", X"0c", X"ed", X"ad", X"6a", 
    X"ae", X"6b", X"8d", X"03", X"8e", X"04", X"1d", X"bd", 
    X"ff", X"01", X"1e", X"eb", X"4c", X"70", X"03", X"02", 
    X"0c", X"ed", X"75", X"82", X"20", X"c0", X"06", X"c0", 
    X"05", X"12", X"0c", X"3b", X"d0", X"05", X"d0", X"06", 
    X"80", X"e0", X"8f", X"82", X"12", X"0c", X"3b", X"02", 
    X"0c", X"ed", X"85", X"4e", X"82", X"85", X"4f", X"83", 
    X"22", X"aa", X"82", X"ab", X"83", X"12", X"14", X"d9", 
    X"60", X"03", X"a3", X"80", X"f8", X"c3", X"e5", X"82", 
    X"9a", X"f5", X"82", X"e5", X"83", X"9b", X"f5", X"83", 
    X"22", X"20", X"f7", X"14", X"30", X"f6", X"14", X"88", 
    X"83", X"a8", X"82", X"20", X"f5", X"07", X"e6", X"a8", 
    X"83", X"75", X"83", X"00", X"22", X"e2", X"80", X"f7", 
    X"e4", X"93", X"22", X"e0", X"22", X"75", X"82", X"00", 
    X"22", X"0a", X"00", X"3e", X"20", X"43", X"35", X"32", 
    X"20", X"6f", X"6e", X"20", X"46", X"50", X"47", X"41", 
    X"20", X"70", X"72", X"6f", X"6a", X"65", X"63", X"74", 
    X"20", X"2d", X"2d", X"20", X"46", X"35", X"32", X"30", 
    X"20", X"63", X"6a", X"68", X"0a", X"00", X"3e", X"20", 
    X"76", X"61", X"6c", X"69", X"64", X"20", X"63", X"6f", 
    X"6d", X"6d", X"61", X"6e", X"64", X"73", X"3a", X"20", 
    X"6c", X"65", X"64", X"20", X"3c", X"68", X"65", X"78", 
    X"3e", X"2c", X"20", X"73", X"77", X"2c", X"20", X"73", 
    X"65", X"63", X"6f", X"6e", X"64", X"73", X"2c", X"20", 
    X"0a", X"00", X"3e", X"20", X"76", X"61", X"6c", X"69", 
    X"64", X"20", X"63", X"6f", X"6d", X"6d", X"61", X"6e", 
    X"64", X"73", X"3a", X"20", X"65", X"6e", X"6c", X"63", 
    X"64", X"20", X"3c", X"68", X"65", X"78", X"3e", X"2c", 
    X"20", X"50", X"30", X"20", X"3c", X"68", X"65", X"78", 
    X"3e", X"2c", X"20", X"50", X"31", X"20", X"3c", X"68", 
    X"65", X"78", X"3e", X"0a", X"00", X"3e", X"20", X"72", 
    X"78", X"20", X"3d", X"20", X"30", X"78", X"25", X"30", 
    X"32", X"78", X"20", X"6e", X"75", X"6d", X"20", X"3d", 
    X"20", X"25", X"64", X"0a", X"00", X"20", X"00", X"3e", 
    X"20", X"61", X"72", X"67", X"76", X"5b", X"30", X"5d", 
    X"20", X"3d", X"20", X"25", X"73", X"0a", X"00", X"3e", 
    X"20", X"61", X"72", X"67", X"76", X"5b", X"31", X"5d", 
    X"20", X"3d", X"20", X"25", X"73", X"0a", X"00", X"6c", 
    X"65", X"64", X"00", X"3e", X"20", X"6c", X"65", X"64", 
    X"20", X"3d", X"20", X"25", X"78", X"0a", X"00", X"73", 
    X"77", X"00", X"3e", X"20", X"73", X"77", X"20", X"3d", 
    X"20", X"25", X"78", X"0a", X"00", X"73", X"65", X"63", 
    X"6f", X"6e", X"64", X"73", X"00", X"3e", X"20", X"73", 
    X"65", X"63", X"6f", X"6e", X"64", X"73", X"20", X"3d", 
    X"20", X"25", X"64", X"0a", X"00", X"50", X"30", X"00", 
    X"3e", X"20", X"50", X"30", X"20", X"3d", X"20", X"25", 
    X"64", X"0a", X"00", X"50", X"31", X"00", X"3e", X"20", 
    X"50", X"31", X"20", X"3d", X"20", X"25", X"64", X"0a", 
    X"00", X"65", X"6e", X"6c", X"63", X"64", X"00", X"3e", 
    X"20", X"65", X"6e", X"6c", X"63", X"64", X"20", X"3d", 
    X"20", X"25", X"64", X"0a", X"00", X"3e", X"20", X"62", 
    X"61", X"63", X"6b", X"73", X"70", X"61", X"63", X"65", 
    X"0a", X"00", X"3c", X"4e", X"4f", X"20", X"46", X"4c", 
    X"4f", X"41", X"54", X"3e", X"00" 
);


end package obj_code_pkg;
